module approx_fa_119_0(X, Y, Z, S, Cout);
input X, Y, Z;
output S, Cout;
assign Cout = 0| (~X & ~Y & Z) | (~X & Y & ~Z) | (~X & Y & Z) | (X & ~Y & Z) | (X & Y & ~Z) | (X & Y & Z) ;
assign S = 0 ;
endmodule
//Compilation time: 2020-12-21 20:54:37
//Compilation SHA256 message digest: a3b96163f4df0c250d004b4f2251d595f41e522f2c4c62c3e7bbdda690c221f0
/*----------------------------------------------------------------------------
Copyright (c) 2019-2020 University of Bremen, Germany.
Copyright (c) 2020 Johannes Kepler University Linz, Austria.
This file has been generated with GenMul.
You can find GenMul at: http://www.sca-verification.org/genmul
Contact us at genmul@sca-verification.org

  First input length: 16
  second input length: 16
  Partial product generator: Unsigned simple partial product generator [U_SP]
  Partial product accumulator: Dadda tree [DT]
  Final stage adder: Ripple carry adder [RC]
----------------------------------------------------------------------------*/
module FullAdder(X, Y, Z, S, C);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule



module U_SP_16_16(IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30);
  input [15:0] IN1;
  input [15:0] IN2;
  output [0:0] P0;
  output [1:0] P1;
  output [2:0] P2;
  output [3:0] P3;
  output [4:0] P4;
  output [5:0] P5;
  output [6:0] P6;
  output [7:0] P7;
  output [8:0] P8;
  output [9:0] P9;
  output [10:0] P10;
  output [11:0] P11;
  output [12:0] P12;
  output [13:0] P13;
  output [14:0] P14;
  output [15:0] P15;
  output [14:0] P16;
  output [13:0] P17;
  output [12:0] P18;
  output [11:0] P19;
  output [10:0] P20;
  output [9:0] P21;
  output [8:0] P22;
  output [7:0] P23;
  output [6:0] P24;
  output [5:0] P25;
  output [4:0] P26;
  output [3:0] P27;
  output [2:0] P28;
  output [1:0] P29;
  output [0:0] P30;
  assign P0[0] = IN1[0]&IN2[0];
  assign P1[0] = IN1[0]&IN2[1];
  assign P2[0] = IN1[0]&IN2[2];
  assign P3[0] = IN1[0]&IN2[3];
  assign P4[0] = IN1[0]&IN2[4];
  assign P5[0] = IN1[0]&IN2[5];
  assign P6[0] = IN1[0]&IN2[6];
  assign P7[0] = IN1[0]&IN2[7];
  assign P8[0] = IN1[0]&IN2[8];
  assign P9[0] = IN1[0]&IN2[9];
  assign P10[0] = IN1[0]&IN2[10];
  assign P11[0] = IN1[0]&IN2[11];
  assign P12[0] = IN1[0]&IN2[12];
  assign P13[0] = IN1[0]&IN2[13];
  assign P14[0] = IN1[0]&IN2[14];
  assign P15[0] = IN1[0]&IN2[15];
  assign P1[1] = IN1[1]&IN2[0];
  assign P2[1] = IN1[1]&IN2[1];
  assign P3[1] = IN1[1]&IN2[2];
  assign P4[1] = IN1[1]&IN2[3];
  assign P5[1] = IN1[1]&IN2[4];
  assign P6[1] = IN1[1]&IN2[5];
  assign P7[1] = IN1[1]&IN2[6];
  assign P8[1] = IN1[1]&IN2[7];
  assign P9[1] = IN1[1]&IN2[8];
  assign P10[1] = IN1[1]&IN2[9];
  assign P11[1] = IN1[1]&IN2[10];
  assign P12[1] = IN1[1]&IN2[11];
  assign P13[1] = IN1[1]&IN2[12];
  assign P14[1] = IN1[1]&IN2[13];
  assign P15[1] = IN1[1]&IN2[14];
  assign P16[0] = IN1[1]&IN2[15];
  assign P2[2] = IN1[2]&IN2[0];
  assign P3[2] = IN1[2]&IN2[1];
  assign P4[2] = IN1[2]&IN2[2];
  assign P5[2] = IN1[2]&IN2[3];
  assign P6[2] = IN1[2]&IN2[4];
  assign P7[2] = IN1[2]&IN2[5];
  assign P8[2] = IN1[2]&IN2[6];
  assign P9[2] = IN1[2]&IN2[7];
  assign P10[2] = IN1[2]&IN2[8];
  assign P11[2] = IN1[2]&IN2[9];
  assign P12[2] = IN1[2]&IN2[10];
  assign P13[2] = IN1[2]&IN2[11];
  assign P14[2] = IN1[2]&IN2[12];
  assign P15[2] = IN1[2]&IN2[13];
  assign P16[1] = IN1[2]&IN2[14];
  assign P17[0] = IN1[2]&IN2[15];
  assign P3[3] = IN1[3]&IN2[0];
  assign P4[3] = IN1[3]&IN2[1];
  assign P5[3] = IN1[3]&IN2[2];
  assign P6[3] = IN1[3]&IN2[3];
  assign P7[3] = IN1[3]&IN2[4];
  assign P8[3] = IN1[3]&IN2[5];
  assign P9[3] = IN1[3]&IN2[6];
  assign P10[3] = IN1[3]&IN2[7];
  assign P11[3] = IN1[3]&IN2[8];
  assign P12[3] = IN1[3]&IN2[9];
  assign P13[3] = IN1[3]&IN2[10];
  assign P14[3] = IN1[3]&IN2[11];
  assign P15[3] = IN1[3]&IN2[12];
  assign P16[2] = IN1[3]&IN2[13];
  assign P17[1] = IN1[3]&IN2[14];
  assign P18[0] = IN1[3]&IN2[15];
  assign P4[4] = IN1[4]&IN2[0];
  assign P5[4] = IN1[4]&IN2[1];
  assign P6[4] = IN1[4]&IN2[2];
  assign P7[4] = IN1[4]&IN2[3];
  assign P8[4] = IN1[4]&IN2[4];
  assign P9[4] = IN1[4]&IN2[5];
  assign P10[4] = IN1[4]&IN2[6];
  assign P11[4] = IN1[4]&IN2[7];
  assign P12[4] = IN1[4]&IN2[8];
  assign P13[4] = IN1[4]&IN2[9];
  assign P14[4] = IN1[4]&IN2[10];
  assign P15[4] = IN1[4]&IN2[11];
  assign P16[3] = IN1[4]&IN2[12];
  assign P17[2] = IN1[4]&IN2[13];
  assign P18[1] = IN1[4]&IN2[14];
  assign P19[0] = IN1[4]&IN2[15];
  assign P5[5] = IN1[5]&IN2[0];
  assign P6[5] = IN1[5]&IN2[1];
  assign P7[5] = IN1[5]&IN2[2];
  assign P8[5] = IN1[5]&IN2[3];
  assign P9[5] = IN1[5]&IN2[4];
  assign P10[5] = IN1[5]&IN2[5];
  assign P11[5] = IN1[5]&IN2[6];
  assign P12[5] = IN1[5]&IN2[7];
  assign P13[5] = IN1[5]&IN2[8];
  assign P14[5] = IN1[5]&IN2[9];
  assign P15[5] = IN1[5]&IN2[10];
  assign P16[4] = IN1[5]&IN2[11];
  assign P17[3] = IN1[5]&IN2[12];
  assign P18[2] = IN1[5]&IN2[13];
  assign P19[1] = IN1[5]&IN2[14];
  assign P20[0] = IN1[5]&IN2[15];
  assign P6[6] = IN1[6]&IN2[0];
  assign P7[6] = IN1[6]&IN2[1];
  assign P8[6] = IN1[6]&IN2[2];
  assign P9[6] = IN1[6]&IN2[3];
  assign P10[6] = IN1[6]&IN2[4];
  assign P11[6] = IN1[6]&IN2[5];
  assign P12[6] = IN1[6]&IN2[6];
  assign P13[6] = IN1[6]&IN2[7];
  assign P14[6] = IN1[6]&IN2[8];
  assign P15[6] = IN1[6]&IN2[9];
  assign P16[5] = IN1[6]&IN2[10];
  assign P17[4] = IN1[6]&IN2[11];
  assign P18[3] = IN1[6]&IN2[12];
  assign P19[2] = IN1[6]&IN2[13];
  assign P20[1] = IN1[6]&IN2[14];
  assign P21[0] = IN1[6]&IN2[15];
  assign P7[7] = IN1[7]&IN2[0];
  assign P8[7] = IN1[7]&IN2[1];
  assign P9[7] = IN1[7]&IN2[2];
  assign P10[7] = IN1[7]&IN2[3];
  assign P11[7] = IN1[7]&IN2[4];
  assign P12[7] = IN1[7]&IN2[5];
  assign P13[7] = IN1[7]&IN2[6];
  assign P14[7] = IN1[7]&IN2[7];
  assign P15[7] = IN1[7]&IN2[8];
  assign P16[6] = IN1[7]&IN2[9];
  assign P17[5] = IN1[7]&IN2[10];
  assign P18[4] = IN1[7]&IN2[11];
  assign P19[3] = IN1[7]&IN2[12];
  assign P20[2] = IN1[7]&IN2[13];
  assign P21[1] = IN1[7]&IN2[14];
  assign P22[0] = IN1[7]&IN2[15];
  assign P8[8] = IN1[8]&IN2[0];
  assign P9[8] = IN1[8]&IN2[1];
  assign P10[8] = IN1[8]&IN2[2];
  assign P11[8] = IN1[8]&IN2[3];
  assign P12[8] = IN1[8]&IN2[4];
  assign P13[8] = IN1[8]&IN2[5];
  assign P14[8] = IN1[8]&IN2[6];
  assign P15[8] = IN1[8]&IN2[7];
  assign P16[7] = IN1[8]&IN2[8];
  assign P17[6] = IN1[8]&IN2[9];
  assign P18[5] = IN1[8]&IN2[10];
  assign P19[4] = IN1[8]&IN2[11];
  assign P20[3] = IN1[8]&IN2[12];
  assign P21[2] = IN1[8]&IN2[13];
  assign P22[1] = IN1[8]&IN2[14];
  assign P23[0] = IN1[8]&IN2[15];
  assign P9[9] = IN1[9]&IN2[0];
  assign P10[9] = IN1[9]&IN2[1];
  assign P11[9] = IN1[9]&IN2[2];
  assign P12[9] = IN1[9]&IN2[3];
  assign P13[9] = IN1[9]&IN2[4];
  assign P14[9] = IN1[9]&IN2[5];
  assign P15[9] = IN1[9]&IN2[6];
  assign P16[8] = IN1[9]&IN2[7];
  assign P17[7] = IN1[9]&IN2[8];
  assign P18[6] = IN1[9]&IN2[9];
  assign P19[5] = IN1[9]&IN2[10];
  assign P20[4] = IN1[9]&IN2[11];
  assign P21[3] = IN1[9]&IN2[12];
  assign P22[2] = IN1[9]&IN2[13];
  assign P23[1] = IN1[9]&IN2[14];
  assign P24[0] = IN1[9]&IN2[15];
  assign P10[10] = IN1[10]&IN2[0];
  assign P11[10] = IN1[10]&IN2[1];
  assign P12[10] = IN1[10]&IN2[2];
  assign P13[10] = IN1[10]&IN2[3];
  assign P14[10] = IN1[10]&IN2[4];
  assign P15[10] = IN1[10]&IN2[5];
  assign P16[9] = IN1[10]&IN2[6];
  assign P17[8] = IN1[10]&IN2[7];
  assign P18[7] = IN1[10]&IN2[8];
  assign P19[6] = IN1[10]&IN2[9];
  assign P20[5] = IN1[10]&IN2[10];
  assign P21[4] = IN1[10]&IN2[11];
  assign P22[3] = IN1[10]&IN2[12];
  assign P23[2] = IN1[10]&IN2[13];
  assign P24[1] = IN1[10]&IN2[14];
  assign P25[0] = IN1[10]&IN2[15];
  assign P11[11] = IN1[11]&IN2[0];
  assign P12[11] = IN1[11]&IN2[1];
  assign P13[11] = IN1[11]&IN2[2];
  assign P14[11] = IN1[11]&IN2[3];
  assign P15[11] = IN1[11]&IN2[4];
  assign P16[10] = IN1[11]&IN2[5];
  assign P17[9] = IN1[11]&IN2[6];
  assign P18[8] = IN1[11]&IN2[7];
  assign P19[7] = IN1[11]&IN2[8];
  assign P20[6] = IN1[11]&IN2[9];
  assign P21[5] = IN1[11]&IN2[10];
  assign P22[4] = IN1[11]&IN2[11];
  assign P23[3] = IN1[11]&IN2[12];
  assign P24[2] = IN1[11]&IN2[13];
  assign P25[1] = IN1[11]&IN2[14];
  assign P26[0] = IN1[11]&IN2[15];
  assign P12[12] = IN1[12]&IN2[0];
  assign P13[12] = IN1[12]&IN2[1];
  assign P14[12] = IN1[12]&IN2[2];
  assign P15[12] = IN1[12]&IN2[3];
  assign P16[11] = IN1[12]&IN2[4];
  assign P17[10] = IN1[12]&IN2[5];
  assign P18[9] = IN1[12]&IN2[6];
  assign P19[8] = IN1[12]&IN2[7];
  assign P20[7] = IN1[12]&IN2[8];
  assign P21[6] = IN1[12]&IN2[9];
  assign P22[5] = IN1[12]&IN2[10];
  assign P23[4] = IN1[12]&IN2[11];
  assign P24[3] = IN1[12]&IN2[12];
  assign P25[2] = IN1[12]&IN2[13];
  assign P26[1] = IN1[12]&IN2[14];
  assign P27[0] = IN1[12]&IN2[15];
  assign P13[13] = IN1[13]&IN2[0];
  assign P14[13] = IN1[13]&IN2[1];
  assign P15[13] = IN1[13]&IN2[2];
  assign P16[12] = IN1[13]&IN2[3];
  assign P17[11] = IN1[13]&IN2[4];
  assign P18[10] = IN1[13]&IN2[5];
  assign P19[9] = IN1[13]&IN2[6];
  assign P20[8] = IN1[13]&IN2[7];
  assign P21[7] = IN1[13]&IN2[8];
  assign P22[6] = IN1[13]&IN2[9];
  assign P23[5] = IN1[13]&IN2[10];
  assign P24[4] = IN1[13]&IN2[11];
  assign P25[3] = IN1[13]&IN2[12];
  assign P26[2] = IN1[13]&IN2[13];
  assign P27[1] = IN1[13]&IN2[14];
  assign P28[0] = IN1[13]&IN2[15];
  assign P14[14] = IN1[14]&IN2[0];
  assign P15[14] = IN1[14]&IN2[1];
  assign P16[13] = IN1[14]&IN2[2];
  assign P17[12] = IN1[14]&IN2[3];
  assign P18[11] = IN1[14]&IN2[4];
  assign P19[10] = IN1[14]&IN2[5];
  assign P20[9] = IN1[14]&IN2[6];
  assign P21[8] = IN1[14]&IN2[7];
  assign P22[7] = IN1[14]&IN2[8];
  assign P23[6] = IN1[14]&IN2[9];
  assign P24[5] = IN1[14]&IN2[10];
  assign P25[4] = IN1[14]&IN2[11];
  assign P26[3] = IN1[14]&IN2[12];
  assign P27[2] = IN1[14]&IN2[13];
  assign P28[1] = IN1[14]&IN2[14];
  assign P29[0] = IN1[14]&IN2[15];
  assign P15[15] = IN1[15]&IN2[0];
  assign P16[14] = IN1[15]&IN2[1];
  assign P17[13] = IN1[15]&IN2[2];
  assign P18[12] = IN1[15]&IN2[3];
  assign P19[11] = IN1[15]&IN2[4];
  assign P20[10] = IN1[15]&IN2[5];
  assign P21[9] = IN1[15]&IN2[6];
  assign P22[8] = IN1[15]&IN2[7];
  assign P23[7] = IN1[15]&IN2[8];
  assign P24[6] = IN1[15]&IN2[9];
  assign P25[5] = IN1[15]&IN2[10];
  assign P26[4] = IN1[15]&IN2[11];
  assign P27[3] = IN1[15]&IN2[12];
  assign P28[2] = IN1[15]&IN2[13];
  assign P29[1] = IN1[15]&IN2[14];
  assign P30[0] = IN1[15]&IN2[15];

endmodule
module DT(IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, IN8, IN9, IN10, IN11, IN12, IN13, IN14, IN15, IN16, IN17, IN18, IN19, IN20, IN21, IN22, IN23, IN24, IN25, IN26, IN27, IN28, IN29, IN30, Out1, Out2);
  input [0:0] IN0;
  input [1:0] IN1;
  input [2:0] IN2;
  input [3:0] IN3;
  input [4:0] IN4;
  input [5:0] IN5;
  input [6:0] IN6;
  input [7:0] IN7;
  input [8:0] IN8;
  input [9:0] IN9;
  input [10:0] IN10;
  input [11:0] IN11;
  input [12:0] IN12;
  input [13:0] IN13;
  input [14:0] IN14;
  input [15:0] IN15;
  input [14:0] IN16;
  input [13:0] IN17;
  input [12:0] IN18;
  input [11:0] IN19;
  input [10:0] IN20;
  input [9:0] IN21;
  input [8:0] IN22;
  input [7:0] IN23;
  input [6:0] IN24;
  input [5:0] IN25;
  input [4:0] IN26;
  input [3:0] IN27;
  input [2:0] IN28;
  input [1:0] IN29;
  input [0:0] IN30;
  output [30:0] Out1;
  output [29:0] Out2;
  wire w256;
  wire w257;
  wire w258;
  wire w259;
  wire w260;
  wire w261;
  wire w262;
  wire w263;
  wire w264;
  wire w265;
  wire w266;
  wire w267;
  wire w268;
  wire w269;
  wire w270;
  wire w271;
  wire w272;
  wire w273;
  wire w274;
  wire w275;
  wire w276;
  wire w277;
  wire w278;
  wire w279;
  wire w280;
  wire w281;
  wire w282;
  wire w283;
  wire w284;
  wire w285;
  wire w286;
  wire w287;
  wire w288;
  wire w289;
  wire w290;
  wire w291;
  wire w292;
  wire w293;
  wire w294;
  wire w295;
  wire w296;
  wire w297;
  wire w298;
  wire w299;
  wire w300;
  wire w301;
  wire w302;
  wire w303;
  wire w304;
  wire w305;
  wire w306;
  wire w307;
  wire w308;
  wire w309;
  wire w310;
  wire w311;
  wire w312;
  wire w313;
  wire w314;
  wire w315;
  wire w316;
  wire w317;
  wire w318;
  wire w319;
  wire w320;
  wire w321;
  wire w322;
  wire w323;
  wire w324;
  wire w325;
  wire w326;
  wire w327;
  wire w328;
  wire w329;
  wire w330;
  wire w331;
  wire w332;
  wire w333;
  wire w334;
  wire w335;
  wire w336;
  wire w337;
  wire w338;
  wire w339;
  wire w340;
  wire w341;
  wire w342;
  wire w343;
  wire w344;
  wire w345;
  wire w346;
  wire w347;
  wire w348;
  wire w349;
  wire w350;
  wire w351;
  wire w352;
  wire w353;
  wire w354;
  wire w355;
  wire w356;
  wire w357;
  wire w358;
  wire w359;
  wire w360;
  wire w361;
  wire w362;
  wire w363;
  wire w364;
  wire w365;
  wire w366;
  wire w367;
  wire w368;
  wire w369;
  wire w370;
  wire w371;
  wire w372;
  wire w373;
  wire w374;
  wire w375;
  wire w376;
  wire w377;
  wire w378;
  wire w379;
  wire w380;
  wire w381;
  wire w382;
  wire w383;
  wire w384;
  wire w385;
  wire w386;
  wire w387;
  wire w388;
  wire w389;
  wire w390;
  wire w391;
  wire w392;
  wire w393;
  wire w394;
  wire w395;
  wire w396;
  wire w397;
  wire w398;
  wire w399;
  wire w400;
  wire w401;
  wire w402;
  wire w403;
  wire w404;
  wire w405;
  wire w406;
  wire w407;
  wire w408;
  wire w409;
  wire w410;
  wire w411;
  wire w412;
  wire w413;
  wire w414;
  wire w415;
  wire w416;
  wire w417;
  wire w418;
  wire w419;
  wire w420;
  wire w421;
  wire w422;
  wire w423;
  wire w424;
  wire w425;
  wire w426;
  wire w427;
  wire w428;
  wire w429;
  wire w430;
  wire w431;
  wire w432;
  wire w433;
  wire w434;
  wire w435;
  wire w436;
  wire w437;
  wire w438;
  wire w439;
  wire w440;
  wire w441;
  wire w442;
  wire w443;
  wire w444;
  wire w445;
  wire w446;
  wire w447;
  wire w448;
  wire w449;
  wire w450;
  wire w451;
  wire w452;
  wire w453;
  wire w454;
  wire w455;
  wire w456;
  wire w457;
  wire w458;
  wire w459;
  wire w460;
  wire w461;
  wire w462;
  wire w463;
  wire w464;
  wire w465;
  wire w466;
  wire w467;
  wire w468;
  wire w469;
  wire w470;
  wire w471;
  wire w472;
  wire w473;
  wire w474;
  wire w475;
  wire w476;
  wire w477;
  wire w478;
  wire w479;
  wire w480;
  wire w481;
  wire w482;
  wire w483;
  wire w484;
  wire w485;
  wire w486;
  wire w487;
  wire w488;
  wire w489;
  wire w490;
  wire w491;
  wire w492;
  wire w493;
  wire w494;
  wire w495;
  wire w496;
  wire w497;
  wire w498;
  wire w499;
  wire w500;
  wire w501;
  wire w502;
  wire w503;
  wire w504;
  wire w505;
  wire w506;
  wire w507;
  wire w508;
  wire w509;
  wire w510;
  wire w511;
  wire w512;
  wire w513;
  wire w514;
  wire w515;
  wire w516;
  wire w517;
  wire w518;
  wire w519;
  wire w520;
  wire w521;
  wire w522;
  wire w523;
  wire w524;
  wire w525;
  wire w526;
  wire w527;
  wire w528;
  wire w529;
  wire w530;
  wire w531;
  wire w532;
  wire w533;
  wire w534;
  wire w535;
  wire w536;
  wire w537;
  wire w538;
  wire w539;
  wire w540;
  wire w541;
  wire w542;
  wire w543;
  wire w544;
  wire w545;
  wire w546;
  wire w547;
  wire w548;
  wire w549;
  wire w550;
  wire w551;
  wire w552;
  wire w553;
  wire w554;
  wire w555;
  wire w556;
  wire w557;
  wire w558;
  wire w559;
  wire w560;
  wire w561;
  wire w562;
  wire w563;
  wire w564;
  wire w565;
  wire w566;
  wire w567;
  wire w568;
  wire w569;
  wire w570;
  wire w571;
  wire w572;
  wire w573;
  wire w574;
  wire w575;
  wire w576;
  wire w577;
  wire w578;
  wire w579;
  wire w580;
  wire w581;
  wire w582;
  wire w583;
  wire w584;
  wire w585;
  wire w586;
  wire w587;
  wire w588;
  wire w589;
  wire w590;
  wire w591;
  wire w592;
  wire w593;
  wire w594;
  wire w595;
  wire w596;
  wire w597;
  wire w598;
  wire w599;
  wire w600;
  wire w601;
  wire w602;
  wire w603;
  wire w604;
  wire w605;
  wire w606;
  wire w607;
  wire w608;
  wire w609;
  wire w610;
  wire w611;
  wire w612;
  wire w613;
  wire w614;
  wire w615;
  wire w616;
  wire w617;
  wire w618;
  wire w619;

  // STAGE 1 
  approx_fa_119_0 L13S1A1 (IN13[0], IN13[1], 1'b0, w256, w257);
  approx_fa_119_0 L14S1A1 (IN14[0], IN14[1], IN14[2], w258, w259);
  approx_fa_119_0 L14S1A2 (IN14[3], IN14[4], 1'b0, w260, w261);
  approx_fa_119_0 L15S1A1 (IN15[0], IN15[1], IN15[2], w262, w263);
  approx_fa_119_0 L15S1A2 (IN15[3], IN15[4], IN15[5], w264, w265);
  approx_fa_119_0 L15S1A3 (IN15[6], IN15[7], 1'b0, w266, w267);
  approx_fa_119_0 L16S1A1 (IN16[0], IN16[1], IN16[2], w268, w269);
  approx_fa_119_0 L16S1A2 (IN16[3], IN16[4], IN16[5], w270, w271);
  approx_fa_119_0 L16S1A3 (IN16[6], IN16[7], 1'b0, w272, w273);
  approx_fa_119_0 L17S1A1 (IN17[0], IN17[1], IN17[2], w274, w275);
  approx_fa_119_0 L17S1A2 (IN17[3], IN17[4], IN17[5], w276, w277);
  approx_fa_119_0 L18S1A1 (IN18[0], IN18[1], IN18[2], w278, w279);

  // STAGE 2 
  approx_fa_119_0 L9S2A1 (IN9[0], IN9[1], 1'b0, w280, w281);
  approx_fa_119_0 L10S2A1 (IN10[0], IN10[1], IN10[2], w282, w283);
  approx_fa_119_0 L10S2A2 (IN10[3], IN10[4], 1'b0, w284, w285);
  approx_fa_119_0 L11S2A1 (IN11[0], IN11[1], IN11[2], w286, w287);
  approx_fa_119_0 L11S2A2 (IN11[3], IN11[4], IN11[5], w288, w289);
  approx_fa_119_0 L11S2A3 (IN11[6], IN11[7], 1'b0, w290, w291);
  approx_fa_119_0 L12S2A1 (IN12[0], IN12[1], IN12[2], w292, w293);
  approx_fa_119_0 L12S2A2 (IN12[3], IN12[4], IN12[5], w294, w295);
  approx_fa_119_0 L12S2A3 (IN12[6], IN12[7], IN12[8], w296, w297);
  approx_fa_119_0 L12S2A4 (IN12[9], IN12[10], 1'b0, w298, w299);
  approx_fa_119_0 L13S2A1 (IN13[2], IN13[3], IN13[4], w300, w301);
  approx_fa_119_0 L13S2A2 (IN13[5], IN13[6], IN13[7], w302, w303);
  approx_fa_119_0 L13S2A3 (IN13[8], IN13[9], IN13[10], w304, w305);
  approx_fa_119_0 L13S2A4 (IN13[11], IN13[12], IN13[13], w306, w307);
  approx_fa_119_0 L14S2A1 (IN14[5], IN14[6], IN14[7], w308, w309);
  approx_fa_119_0 L14S2A2 (IN14[8], IN14[9], IN14[10], w310, w311);
  approx_fa_119_0 L14S2A3 (IN14[11], IN14[12], IN14[13], w312, w313);
  approx_fa_119_0 L14S2A4 (IN14[14], w257, w258, w314, w315);
  approx_fa_119_0 L15S2A1 (IN15[8], IN15[9], IN15[10], w316, w317);
  approx_fa_119_0 L15S2A2 (IN15[11], IN15[12], IN15[13], w318, w319);
  approx_fa_119_0 L15S2A3 (IN15[14], IN15[15], w259, w320, w321);
  approx_fa_119_0 L15S2A4 (w261, w262, w264, w322, w323);
  approx_fa_119_0 L16S2A1 (IN16[8], IN16[9], IN16[10], w324, w325);
  approx_fa_119_0 L16S2A2 (IN16[11], IN16[12], IN16[13], w326, w327);
  approx_fa_119_0 L16S2A3 (IN16[14], w263, w265, w328, w329);
  approx_fa_119_0 L16S2A4 (w267, w268, w270, w330, w331);
  approx_fa_119_0 L17S2A1 (IN17[6], IN17[7], IN17[8], w332, w333);
  approx_fa_119_0 L17S2A2 (IN17[9], IN17[10], IN17[11], w334, w335);
  approx_fa_119_0 L17S2A3 (IN17[12], IN17[13], w269, w336, w337);
  approx_fa_119_0 L17S2A4 (w271, w273, w274, w338, w339);
  approx_fa_119_0 L18S2A1 (IN18[3], IN18[4], IN18[5], w340, w341);
  approx_fa_119_0 L18S2A2 (IN18[6], IN18[7], IN18[8], w342, w343);
  approx_fa_119_0 L18S2A3 (IN18[9], IN18[10], IN18[11], w344, w345);
  approx_fa_119_0 L18S2A4 (IN18[12], w275, w277, w346, w347);
  approx_fa_119_0 L19S2A1 (IN19[0], IN19[1], IN19[2], w348, w349);
  approx_fa_119_0 L19S2A2 (IN19[3], IN19[4], IN19[5], w350, w351);
  approx_fa_119_0 L19S2A3 (IN19[6], IN19[7], IN19[8], w352, w353);
  approx_fa_119_0 L19S2A4 (IN19[9], IN19[10], IN19[11], w354, w355);
  approx_fa_119_0 L20S2A1 (IN20[0], IN20[1], IN20[2], w356, w357);
  approx_fa_119_0 L20S2A2 (IN20[3], IN20[4], IN20[5], w358, w359);
  approx_fa_119_0 L20S2A3 (IN20[6], IN20[7], IN20[8], w360, w361);
  FullAdder L21S2A1 (IN21[0], IN21[1], IN21[2], w362, w363);
  FullAdder L21S2A2 (IN21[3], IN21[4], IN21[5], w364, w365);
  FullAdder L22S2A1 (IN22[0], IN22[1], IN22[2], w366, w367);

  // STAGE 3
  approx_fa_119_0 L6S3A1 (IN6[0], IN6[1], 1'b0, w368, w369);
  approx_fa_119_0 L7S3A1 (IN7[0], IN7[1], IN7[2], w370, w371);
  approx_fa_119_0 L7S3A2 (IN7[3], IN7[4], 1'b0, w372, w373);
  approx_fa_119_0 L8S3A1 (IN8[0], IN8[1], IN8[2], w374, w375);
  approx_fa_119_0 L8S3A2 (IN8[3], IN8[4], IN8[5], w376, w377);
  approx_fa_119_0 L8S3A3 (IN8[6], IN8[7], 1'b0, w378, w379);
  approx_fa_119_0 L9S3A1 (IN9[2], IN9[3], IN9[4], w380, w381);
  approx_fa_119_0 L9S3A2 (IN9[5], IN9[6], IN9[7], w382, w383);
  approx_fa_119_0 L9S3A3 (IN9[8], IN9[9], w280, w384, w385);
  approx_fa_119_0 L10S3A1 (IN10[5], IN10[6], IN10[7], w386, w387);
  approx_fa_119_0 L10S3A2 (IN10[8], IN10[9], IN10[10], w388, w389);
  approx_fa_119_0 L10S3A3 (w281, w282, w284, w390, w391);
  approx_fa_119_0 L11S3A1 (IN11[8], IN11[9], IN11[10], w392, w393);
  approx_fa_119_0 L11S3A2 (IN11[11], w283, w285, w394, w395);
  approx_fa_119_0 L11S3A3 (w286, w288, w290, w396, w397);
  approx_fa_119_0 L12S3A1 (IN12[11], IN12[12], w287, w398, w399);
  approx_fa_119_0 L12S3A2 (w289, w291, w292, w400, w401);
  approx_fa_119_0 L12S3A3 (w294, w296, w298, w402, w403);
  approx_fa_119_0 L13S3A1 (w256, w293, w295, w404, w405);
  approx_fa_119_0 L13S3A2 (w297, w299, w300, w406, w407);
  approx_fa_119_0 L13S3A3 (w302, w304, w306, w408, w409);
  approx_fa_119_0 L14S3A1 (w260, w301, w303, w410, w411);
  approx_fa_119_0 L14S3A2 (w305, w307, w308, w412, w413);
  approx_fa_119_0 L14S3A3 (w310, w312, w314, w414, w415);
  approx_fa_119_0 L15S3A1 (w266, w309, w311, w416, w417);
  approx_fa_119_0 L15S3A2 (w313, w315, w316, w418, w419);
  approx_fa_119_0 L15S3A3 (w318, w320, w322, w420, w421);
  approx_fa_119_0 L16S3A1 (w272, w317, w319, w422, w423);
  approx_fa_119_0 L16S3A2 (w321, w323, w324, w424, w425);
  approx_fa_119_0 L16S3A3 (w326, w328, w330, w426, w427);
  approx_fa_119_0 L17S3A1 (w276, w325, w327, w428, w429);
  approx_fa_119_0 L17S3A2 (w329, w331, w332, w430, w431);
  approx_fa_119_0 L17S3A3 (w334, w336, w338, w432, w433);
  approx_fa_119_0 L18S3A1 (w278, w333, w335, w434, w435);
  approx_fa_119_0 L18S3A2 (w337, w339, w340, w436, w437);
  approx_fa_119_0 L18S3A3 (w342, w344, w346, w438, w439);
  approx_fa_119_0 L19S3A1 (w279, w341, w343, w440, w441);
  approx_fa_119_0 L19S3A2 (w345, w347, w348, w442, w443);
  approx_fa_119_0 L19S3A3 (w350, w352, w354, w444, w445);
  approx_fa_119_0 L20S3A1 (IN20[9], IN20[10], w349, w446, w447);
  approx_fa_119_0 L20S3A2 (w351, w353, w355, w448, w449);
  approx_fa_119_0 L20S3A3 (w356, w358, w360, w450, w451);
  FullAdder L21S3A1 (IN21[6], IN21[7], IN21[8], w452, w453);
  FullAdder L21S3A2 (IN21[9], w357, w359, w454, w455);
  FullAdder L21S3A3 (w361, w362, w364, w456, w457);
  FullAdder L22S3A1 (IN22[3], IN22[4], IN22[5], w458, w459);
  FullAdder L22S3A2 (IN22[6], IN22[7], IN22[8], w460, w461);
  FullAdder L22S3A3 (w363, w365, w366, w462, w463);
  FullAdder L23S3A1 (IN23[0], IN23[1], IN23[2], w464, w465);
  FullAdder L23S3A2 (IN23[3], IN23[4], IN23[5], w466, w467);
  FullAdder L23S3A3 (IN23[6], IN23[7], w367, w468, w469);
  FullAdder L24S3A1 (IN24[0], IN24[1], IN24[2], w470, w471);
  FullAdder L24S3A2 (IN24[3], IN24[4], IN24[5], w472, w473);
  FullAdder L25S3A1 (IN25[0], IN25[1], IN25[2], w474, w475);
  
  // STAGE 4 
  approx_fa_119_0 L4S4A1 (IN4[0], IN4[1], 1'b0, w476, w477);
  approx_fa_119_0 L5S4A1 (IN5[0], IN5[1], IN5[2], w478, w479);
  approx_fa_119_0 L5S4A2 (IN5[3], IN5[4], 1'b0, w480, w481);
  approx_fa_119_0 L6S4A1 (IN6[2], IN6[3], IN6[4], w482, w483);
  approx_fa_119_0 L6S4A2 (IN6[5], IN6[6], w368, w484, w485);
  approx_fa_119_0 L7S4A1 (IN7[5], IN7[6], IN7[7], w486, w487);
  approx_fa_119_0 L7S4A2 (w369, w370, w372, w488, w489);
  approx_fa_119_0 L8S4A1 (IN8[8], w371, w373, w490, w491);
  approx_fa_119_0 L8S4A2 (w374, w376, w378, w492, w493);
  approx_fa_119_0 L9S4A1 (w375, w377, w379, w494, w495);
  approx_fa_119_0 L9S4A2 (w380, w382, w384, w496, w497);
  approx_fa_119_0 L10S4A1 (w381, w383, w385, w498, w499);
  approx_fa_119_0 L10S4A2 (w386, w388, w390, w500, w501);
  approx_fa_119_0 L11S4A1 (w387, w389, w391, w502, w503);
  approx_fa_119_0 L11S4A2 (w392, w394, w396, w504, w505);
  approx_fa_119_0 L12S4A1 (w393, w395, w397, w506, w507);
  approx_fa_119_0 L12S4A2 (w398, w400, w402, w508, w509);
  approx_fa_119_0 L13S4A1 (w399, w401, w403, w510, w511);
  approx_fa_119_0 L13S4A2 (w404, w406, w408, w512, w513);
  approx_fa_119_0 L14S4A1 (w405, w407, w409, w514, w515);
  approx_fa_119_0 L14S4A2 (w410, w412, w414, w516, w517);
  approx_fa_119_0 L15S4A1 (w411, w413, w415, w518, w519);
  approx_fa_119_0 L15S4A2 (w416, w418, w420, w520, w521);
  approx_fa_119_0 L16S4A1 (w417, w419, w421, w522, w523);
  approx_fa_119_0 L16S4A2 (w422, w424, w426, w524, w525);
  approx_fa_119_0 L17S4A1 (w423, w425, w427, w526, w527);
  approx_fa_119_0 L17S4A2 (w428, w430, w432, w528, w529);
  approx_fa_119_0 L18S4A1 (w429, w431, w433, w530, w531);
  approx_fa_119_0 L18S4A2 (w434, w436, w438, w532, w533);
  approx_fa_119_0 L19S4A1 (w435, w437, w439, w534, w535);
  approx_fa_119_0 L19S4A2 (w440, w442, w444, w536, w537);
  approx_fa_119_0 L20S4A1 (w441, w443, w445, w538, w539);
  approx_fa_119_0 L20S4A2 (w446, w448, w450, w540, w541);
  FullAdder L21S4A1 (w447, w449, w451, w542, w543);
  FullAdder L21S4A2 (w452, w454, w456, w544, w545);
  FullAdder L22S4A1 (w453, w455, w457, w546, w547);
  FullAdder L22S4A2 (w458, w460, w462, w548, w549);
  FullAdder L23S4A1 (w459, w461, w463, w550, w551);
  FullAdder L23S4A2 (w464, w466, w468, w552, w553);
  FullAdder L24S4A1 (IN24[6], w465, w467, w554, w555);
  FullAdder L24S4A2 (w469, w470, w472, w556, w557);
  FullAdder L25S4A1 (IN25[3], IN25[4], IN25[5], w558, w559);
  FullAdder L25S4A2 (w471, w473, w474, w560, w561);
  FullAdder L26S4A1 (IN26[0], IN26[1], IN26[2], w562, w563);
  FullAdder L26S4A2 (IN26[3], IN26[4], w475, w564, w565);
  FullAdder L27S4A1 (IN27[0], IN27[1], IN27[2], w566, w567);
 
  // STAGE 5
  approx_fa_119_0 L3S5A1 (IN3[0], IN3[1], 1'b0, w568, w569);
  approx_fa_119_0 L4S5A1 (IN4[2], IN4[3], IN4[4], w570, w571);
  approx_fa_119_0 L5S5A1 (IN5[5], w477, w478, w572, w573);
  approx_fa_119_0 L6S5A1 (w479, w481, w482, w574, w575);
  approx_fa_119_0 L7S5A1 (w483, w485, w486, w576, w577);
  approx_fa_119_0 L8S5A1 (w487, w489, w490, w578, w579);
  approx_fa_119_0 L9S5A1 (w491, w493, w494, w580, w581);
  approx_fa_119_0 L10S5A1 (w495, w497, w498, w582, w583);
  approx_fa_119_0 L11S5A1 (w499, w501, w502, w584, w585);
  approx_fa_119_0 L12S5A1 (w503, w505, w506, w586, w587);
  approx_fa_119_0 L13S5A1 (w507, w509, w510, w588, w589);
  approx_fa_119_0 L14S5A1 (w511, w513, w514, w590, w591);
  approx_fa_119_0 L15S5A1 (w515, w517, w518, w592, w593);
  approx_fa_119_0 L16S5A1 (w519, w521, w522, w594, w595);
  approx_fa_119_0 L17S5A1 (w523, w525, w526, w596, w597);
  approx_fa_119_0 L18S5A1 (w527, w529, w530, w598, w599);
  approx_fa_119_0 L19S5A1 (w531, w533, w534, w600, w601);
  approx_fa_119_0 L20S5A1 (w535, w537, w538, w602, w603);
  FullAdder L21S5A1 (w539, w541, w542, w604, w605);
  FullAdder L22S5A1 (w543, w545, w546, w606, w607);
  FullAdder L23S5A1 (w547, w549, w550, w608, w609);
  FullAdder L24S5A1 (w551, w553, w554, w610, w611);
  FullAdder L25S5A1 (w555, w557, w558, w612, w613);
  FullAdder L26S5A1 (w559, w561, w562, w614, w615);
  FullAdder L27S5A1 (IN27[3], w563, w565, w616, w617);
  FullAdder L28S5A1 (IN28[0], IN28[1], IN28[2], w618, w619);
  
  //STAGE 6
  approx_fa_119_0 L2S6A1 (IN2[0], IN2[1], 1'b0, Out2[1], Out1[3]);
  approx_fa_119_0 L3S6A1 (IN3[2], IN3[3], w568, Out2[2], Out1[4]);
  approx_fa_119_0 L4S6A1 (w476, w569, w570, Out2[3], Out1[5]);
  approx_fa_119_0 L5S6A1 (w480, w571, w572, Out2[4], Out1[6]);
  approx_fa_119_0 L6S6A1 (w484, w573, w574, Out2[5], Out1[7]);
  approx_fa_119_0 L7S6A1 (w488, w575, w576, Out2[6], Out1[8]);
  approx_fa_119_0 L8S6A1 (w492, w577, w578, Out2[7], Out1[9]);
  approx_fa_119_0 L9S6A1 (w496, w579, w580, Out2[8], Out1[10]);
  approx_fa_119_0 L10S6A1 (w500, w581, w582, Out2[9], Out1[11]);
  approx_fa_119_0 L11S6A1 (w504, w583, w584, Out2[10], Out1[12]);
  approx_fa_119_0 L12S6A1 (w508, w585, w586, Out2[11], Out1[13]);
  approx_fa_119_0 L13S6A1 (w512, w587, w588, Out2[12], Out1[14]);
  approx_fa_119_0 L14S6A1 (w516, w589, w590, Out2[13], Out1[15]);
  approx_fa_119_0 L15S6A1 (w520, w591, w592, Out2[14], Out1[16]);
  approx_fa_119_0 L16S6A1 (w524, w593, w594, Out2[15], Out1[17]);
  approx_fa_119_0 L17S6A1 (w528, w595, w596, Out2[16], Out1[18]);
  approx_fa_119_0 L18S6A1 (w532, w597, w598, Out2[17], Out1[19]);
  approx_fa_119_0 L19S6A1 (w536, w599, w600, Out2[18], Out1[20]);
  approx_fa_119_0 L20S6A1 (w540, w601, w602, Out2[19], Out1[21]);
  FullAdder L21S6A1 (w544, w603, w604, Out2[20], Out1[22]);
  FullAdder L22S6A1 (w548, w605, w606, Out2[21], Out1[23]);
  FullAdder L23S6A1 (w552, w607, w608, Out2[22], Out1[24]);
  FullAdder L24S6A1 (w556, w609, w610, Out2[23], Out1[25]);
  FullAdder L25S6A1 (w560, w611, w612, Out2[24], Out1[26]);
  FullAdder L26S6A1 (w564, w613, w614, Out2[25], Out1[27]);
  FullAdder L27S6A1 (w566, w615, w616, Out2[26], Out1[28]);
  FullAdder L28S6A1 (w567, w617, w618, Out2[27], Out1[29]);
  FullAdder L29S6A1 (IN29[0], IN29[1], w619, Out2[28], Out2[29]);
  assign Out1[0] = IN0[0];
  assign Out1[1] = IN1[0];
  assign Out2[0] = IN1[1];
  assign Out1[2] = IN2[2];
  assign Out1[30] = IN30[0];

endmodule
module RC_30_30(IN1, IN2, Out);
  input [29:0] IN1;
  input [29:0] IN2;
  output [30:0] Out;
  wire w61;
  wire w63;
  wire w65;
  wire w67;
  wire w69;
  wire w71;
  wire w73;
  wire w75;
  wire w77;
  wire w79;
  wire w81;
  wire w83;
  wire w85;
  wire w87;
  wire w89;
  wire w91;
  wire w93;
  wire w95;
  wire w97;
  wire w99;
  wire w101;
  wire w103;
  wire w105;
  wire w107;
  wire w109;
  wire w111;
  wire w113;
  wire w115;
  wire w117;
  approx_fa_119_0 L1S7A1 (IN1[0], IN2[0], 1'b0, Out[0], w61);
  approx_fa_119_0 L2S7A1 (IN1[1], IN2[1], w61, Out[1], w63);
  approx_fa_119_0 L3S7A1 (IN1[2], IN2[2], w63, Out[2], w65);
  approx_fa_119_0 L4S7A1 (IN1[3], IN2[3], w65, Out[3], w67);
  approx_fa_119_0 L5S7A1 (IN1[4], IN2[4], w67, Out[4], w69);
  approx_fa_119_0 L6S7A1 (IN1[5], IN2[5], w69, Out[5], w71);
  approx_fa_119_0 L7S7A1 (IN1[6], IN2[6], w71, Out[6], w73);
  approx_fa_119_0 L8S7A1 (IN1[7], IN2[7], w73, Out[7], w75);
  approx_fa_119_0 L9S7A1 (IN1[8], IN2[8], w75, Out[8], w77);
  approx_fa_119_0 L10S7A1 (IN1[9], IN2[9], w77, Out[9], w79);
  approx_fa_119_0 L11S7A1 (IN1[10], IN2[10], w79, Out[10], w81);
  approx_fa_119_0 L12S7A1 (IN1[11], IN2[11], w81, Out[11], w83);
  approx_fa_119_0 L13S7A1 (IN1[12], IN2[12], w83, Out[12], w85);
  approx_fa_119_0 L14S7A1 (IN1[13], IN2[13], w85, Out[13], w87);
  approx_fa_119_0 L15S7A1 (IN1[14], IN2[14], w87, Out[14], w89);
  approx_fa_119_0 L16S7A1 (IN1[15], IN2[15], w89, Out[15], w91);
  approx_fa_119_0 L17S7A1 (IN1[16], IN2[16], w91, Out[16], w93);
  approx_fa_119_0 L18S7A1 (IN1[17], IN2[17], w93, Out[17], w95);
  approx_fa_119_0 L19S7A1 (IN1[18], IN2[18], w95, Out[18], w97);
  approx_fa_119_0 L20S7A1 (IN1[19], IN2[19], w97, Out[19], w99);
  FullAdder L21S7A1 (IN1[20], IN2[20], w99, Out[20], w101);
  FullAdder L22S7A1 (IN1[21], IN2[21], w101, Out[21], w103);
  FullAdder L23S7A1 (IN1[22], IN2[22], w103, Out[22], w105);
  FullAdder L24S7A1 (IN1[23], IN2[23], w105, Out[23], w107);
  FullAdder L25S7A1 (IN1[24], IN2[24], w107, Out[24], w109);
  FullAdder L26S7A1 (IN1[25], IN2[25], w109, Out[25], w111);
  FullAdder L27S7A1 (IN1[26], IN2[26], w111, Out[26], w113);
  FullAdder L28S7A1 (IN1[27], IN2[27], w113, Out[27], w115);
  FullAdder L29S7A1 (IN1[28], IN2[28], w115, Out[28], w117);
  FullAdder L30S7A1 (IN1[29], IN2[29], w117, Out[29], Out[30]);

endmodule
module DT_16_16_20_approx_fa_119_0(IN1, IN2, Out);
  input [15:0] IN1;
  input [15:0] IN2;
  output [31:0] Out;
  wire [0:0] P0;
  wire [1:0] P1;
  wire [2:0] P2;
  wire [3:0] P3;
  wire [4:0] P4;
  wire [5:0] P5;
  wire [6:0] P6;
  wire [7:0] P7;
  wire [8:0] P8;
  wire [9:0] P9;
  wire [10:0] P10;
  wire [11:0] P11;
  wire [12:0] P12;
  wire [13:0] P13;
  wire [14:0] P14;
  wire [15:0] P15;
  wire [14:0] P16;
  wire [13:0] P17;
  wire [12:0] P18;
  wire [11:0] P19;
  wire [10:0] P20;
  wire [9:0] P21;
  wire [8:0] P22;
  wire [7:0] P23;
  wire [6:0] P24;
  wire [5:0] P25;
  wire [4:0] P26;
  wire [3:0] P27;
  wire [2:0] P28;
  wire [1:0] P29;
  wire [0:0] P30;
  wire [30:0] R1;
  wire [29:0] R2;
  wire [31:0] aOut;
  U_SP_16_16 S0 (IN1, IN2 , P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30);
  DT S1 (P0, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, P11, P12, P13, P14, P15, P16, P17, P18, P19, P20, P21, P22, P23, P24, P25, P26, P27, P28, P29, P30, R1, R2);
  RC_30_30 S2 (R1[30:1], R2, aOut[31:1]);
  assign aOut[0] = R1[0];
  assign Out = aOut[31:0];
endmodule

/*---------------------------------------------------------------------------------------------------
This are SHA256 message digests computed for all source files to see the version of a file in genmul.
4164f841dcd2afb1341b584b40f40d82ef4c3d0830615503b45c13f9ff1f0b99 Array.cpp
b66c13355402b785b10523902060ea2b13495e0139581e3e1f9eb511b63091d0 Array.hpp
049f660c454752c510b8d2d7d5474b271804a3f2ef3bbd08b201b27cf5aa953c BrentKungAdder.cpp
542006e2bd9fe43a38fbd454d79c40216e2222968ee81d61ccb8b9f5f7c2cfc0 BrentKungAdder.hpp
dd0e0628729b9c228e1e3e2d8c759e3c5d548b2a7fc7a0ecf965f77c057f8982 CarryLookAhead.cpp
acab3bf6b24f0596013dfce2d21a56d16bc4565d810d7521bef6b645b6192ddf CarryLookAhead.hpp
929ba8b159d43cd1483702c39adf3f3c01a0e029393157d2dff1e576c3784ba2 CarryPredictor.cpp
c674a6131475e399d67794664958ce3992e34ad5a8a276b258f3b65179dbb0d2 CarryPredictor.hpp
7ad1df61ce6dec8970320cdbb0cd1b9d9e1b1aaed8337fad2ba9dc15bebade69 CarrySkipAdder.cpp
ce45d117e5a45c141acb0a305a0a6eaf30ccdc4b387a55bd5ab330672bf3c03a CarrySkipAdder.hpp
227583b37ff516c46466fc5c918ee7605b0476c7e79e1b63b1fc28017046b0d2 CarrySkipAdderVariable.cpp
1812c7c9c45afa80da1317afd4c2210c3583748daed3177e247887653392a938 CarrySkipAdderVariable.hpp
6cb775e3f48c2bc7fe32ff327217939a020f17c5087cc13d0faee3452517d768 component.cpp
209f908d2f1fb45ff2ab578483ac59b4daf3db09b0623e939fe467d8c408a03c component.hpp
1448c3a20470e843c0e3d8e81150aa7ae966b01c0324366ad6d09973635eae33 Dadda.cpp
b409b894cf7e5dd8b1566ad65242d8204a3b10e09218cfdba51d6798420c3db4 Dadda.hpp
e2de7008e12d31cf28e87ddcc91be289718e8c57104720d626d739224e17d237 GenMul.cpp
ca6978e216edf5aa647ec0ac3ce023db92fac8b0514ff9494e53594d0f6870ea GenMul_Emscripten.cpp
59b5e2c157f082415d42add003c3f61c2a59ddcff55d4bce8b87b7769944c265 GenMul_Emscripten.hpp
9f7728b1956d663933ee8c2e36eedbfbf99e183f597155867c1b3ea7b518cfc7 GenMul.hpp
b6c44052471006782baa14f9ee553e9dd2befb5a48caaf3ea08ada0fa333a4b7 KoggeStoneAdder.cpp
39decce3c706b8eafdd039498cb80147312dc279cf9ac722df1d7c5e44ca1eb1 KoggeStoneAdder.hpp
8cd281edd6691072195380d088347b8080c00b9bdc903f9930b6f9b66343a532 LanderFischerAdder.cpp
5a7fd4ccf6aba5d41505bf471d36050ebc082c671b174d26d2afe89d8ab1424f LanderFischerAdder.hpp
e882c7b4ccf415774af64e8554a5d95bc8652feda0a36406f200e95b0228339b main.cpp
bc20681185e8c41a7f23ff828021720d345a078c484211fe91f92bc0bffc69e2 ModuleConnector.cpp
e1e43efd032bbdf2f7cde39e51a5ca384a6f7dbe2bbb2d60b2ce379cba5c5a61 ModuleConnector.hpp
287f82e4c4496d55e1bfa8679ee9e55e472790befa8efd8632594da9f222bcc6 partial.cpp
0f936d14fa3aa23fae3171e401a240bea867f3be47b3cf7302cfabd3cb016a2a partial.hpp
8ce42bf2a0b4a30bf2a9b1371c7e59d94c8b71af34319211923ebc0acae9f0d0 PartialProductGenerator.cpp
0ec3b8793327e4b4e723a90196524386697346d2ab66595de11ae34a7ed16ae2 PartialProductGenerator.hpp
049b30b6e146bee3b19fa21ee9d78e1fba8caf3bf38b0e4a99bc6e35110f8cef PartialProductGeneratorSigned.cpp
b3fd13d4dc90c5708b5905c73a6437578e972e9929a8f5ef40d224277a72b3eb PartialProductGeneratorSigned.hpp
b4d8f357fdd48208ab4dbec18a26d3dd8091c289f388f9bfe66dfe22793c005c RippleCarryAdder.cpp
7a68cc632729d6a10a87e0d6750a3b6bc38ffea3c1adefbb6c04f5c81d6821fd RippleCarryAdder.hpp
02ad7291a8c88d72769d019fcfcb63f20595eeb7f97880174f7080c433adc827 SerialPrefixAdder.cpp
34c8850d96db902dcf9124b07b854739c311e1b984f27ae2cba2c97dac68b528 SerialPrefixAdder.hpp
ce0ae8c29d242e8eda47cc3e9ff06bb052ce1a90f3c8e0cf21ee13c63ddd30e9 VerilogGen.cpp
60865ceaeae304e64ad944fb7b83fda22058c3e042b9e5ad1e2b35effcb79918 VerilogGen.hpp
421854807ffbed49e9450453ff4d7b2fb6cbcff53c1e8cca3299cc3c49d5bb6f Wallace5.cpp
ae5f879f4f6fda292e6394ba3e8df4a50b38d2c1c8f590fbf5752c2109deb398 Wallace5.hpp
53e7bc2a228005f30c0349cd8f1e2f68498141e175ee1c140d3465823cfc44ec Wallace.cpp
f00fd621015cfcf54cda85815dce343d8526c1fee0f7e22a9d98041195b72e1a Wallace.hpp
---------------------------------------------------------------------------------------------------*/

